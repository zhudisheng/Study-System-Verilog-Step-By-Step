module test_operator;
reg [7:0] a,b,c;
initial begin
	a=10;b=11;c=12;
	$display("Assignment Operators:");
	$display("a = 	%d  %d",a,a);
	#10 a += 2;
	$display("a += 	%d  %d",a,a);
	#10 a -= 2;
	$display("a -= 	%d  %d",a,a);
	#10 a *= 2;
	$display("a *= 	%d  %d",a,a);
	#10 a /= 2;
	$display("a /= 	%d  %d",a,a);
	#10 a %= 3;
	$display("a mod= %d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a &= 2;
	$display("a &= 	%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a |= 2;
	$display("a |= 	%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a ^= 2;
	$display("a ^= 	%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a <<= 2;
	$display("a <<=	%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a >>= 2;
	$display("a >>=	%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a <<<= 2;
	$display("a <<<=%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d  %d",a,a);
	#10 a >>>= 2;
	$display("a >>>=%d  %d",a,a);
	#10 a = 'hc3;
	$display("a = 	%d",a);
	$display("a++ :	%d",a++);
	$display("++a :	%d",++a);
	$display("a-- :	%d",a--);
	$display("--a :	%d",--a);
end
endmodule
