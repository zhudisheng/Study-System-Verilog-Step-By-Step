program test;
    initial begin
        $display("hello world!");
    end
endprogram
